* SPICE NETLIST
***************************************

.SUBCKT test_nmos Vout Vd Vg
** N=7 EP=3 IP=0 FDC=1
M0 Vd Vg Vout Vout nch_18_mac L=1.5e-08 W=3.2e-08 $X=2000 $Y=2300 $D=0
.ENDS
***************************************
