* SPICE NETLIST
***************************************

.SUBCKT test_pdio V1 V2
** N=2 EP=2 IP=0 FDC=1
D0 V1 V2 pdio AREA=9e-12 PJ=1.2e-05 $X=780 $Y=-4755 $D=0
.ENDS
***************************************
