* SPICE NETLIST
***************************************

.SUBCKT pnp_CDNS_627487506800 1 2 3
** N=3 EP=3 IP=0 FDC=1
Q0 1 3 2 pnp5 AREA=2.5e-11 $X=2100 $Y=2100 $D=0
.ENDS
***************************************
.SUBCKT test_pnp Vc Vb Ve
** N=3 EP=3 IP=9 FDC=3
X0 Vc Ve Vb pnp_CDNS_627487506800 $T=500 -10700 0 0 $X=500 $Y=-10700
X1 Vc Ve Vb pnp_CDNS_627487506800 $T=10700 -10700 0 0 $X=10700 $Y=-10700
X2 Vc Ve Vb pnp_CDNS_627487506800 $T=20900 -10700 0 0 $X=20900 $Y=-10700
.ENDS
***************************************
